--
-- VHDL Architecture my_project4_lib.controller.b
--
-- Created:
--          by - Wei Guo.UNKNOWN (MSI)
--          at - 17:28:48 03/17/2018
--
-- using Mentor Graphics HDL Designer(TM) 2015.1b (Build 4)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY controller IS
END ENTITY controller;

--
ARCHITECTURE b OF controller IS
BEGIN
END ARCHITECTURE b;

